--
--Written by GowinSynthesis
--Tool Version "V1.9.12 (64-bit)"
--Sun Dec 28 11:45:49 2025

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/SPIMASTER/data/spi_master_top.v"
--file1 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/SPIMASTER/data/spi_master.vp"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
KZTH8QXEnMw1PxgnrUkdNMzkebbM6gz8m9+mugIaCW8/uHKX3Ay/jw/+tZ5wXugrM6q257T0Wwn6
NK5PT4KGfQFYmmpLZpF+A1nIZ3I7Uggr++ZAhhyba/6pEBecmbPG/mfJpPJPkzyxTzpDGOBc1vt6
ogqMVCfBb1cRSautHb2vPBa3JGvPTlhXlx6uCoeMtyoltHfrbtLPodEUVFYJ8V623Sqqu6OkQnvO
CuJOhRyZopKIln4Lkzo8ZKpxIyKbixzGOzt0+nR7XCIv/a7itBtvLCaZzyhN5aCqZftVCn5etR3J
l9Kz4qYcA+9OjInSXp59aTSgCk4qSol+qKkHeQ==

`protect encoding=(enctype="base64", line_length=76, bytes=29840)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
tqapmJUw1+tDb4Xpdo46x6ZjSSLYp3uVEijT+yKmz22zHbOXcwZxdaF6FCFWYAwuS4uhSJCKta6p
7OODehncoswziXANU3GbCl8bgOeuITLQH8glC+zT/Rnpi+7irUA+UBL08h8CrSr9ePIjpkigFHLa
PZoAHKTczZszmDFKoUEWOI3PnJsm+XwYZrTlXM3bRKpKdUmyGm6LWzrBzJpZOm3cINrKYgWCY+t0
k/LKg7FqDkNh/MSVvTNQoS2a7+LKv4uDGjHd0U9LCHXIKwZkhIS9Rd17xxKZ6XQ0jCbFaLAEfH4U
+ipYBfgYDXv/i6MED7nROlNjsmkB3HPX6Di/OB//fhVmnfoe1FNlr89vaofYADlJpS/YECmllrKG
YoenYtznlAFb6eAIZAopmLmw5nBvLpu5RQNEBN2CpCl4G40J50UIetY+99e+taPVNxAfczt6+6GM
e1TLzQH4ZQCDhhJn5D9WomaFQGLmFcVm5cQCAPcFYlHpw3TjOo9kaHLtPjVs7qb2HBBAcnjwo6bC
AxNIADfBgg9ODiH7WMYehzkaLIk1yJGTFpDLD6t827unP5cA+iRB+VVY0I9grZDStzlmu0hhIh4P
0LQZ+FY8Eb21+vPx6yiJslqVt9SjZRuf7Un/9eit+Fv6jSAnzP+k4D3ulg6KVz80zs1ioC7WcTKW
RgsV0Szn1Z/D7IJSP7rDweHUy833Qj0kPYcUH8Xt9FC1wLtyihIftR9ThBpOjj60uGjB6KnzOGbO
m39pPK0NTojPIP73LEMzdsZ/vmB5tLkdSWOu25GlOKHtld2KDvXpQrvug+opFLrdGNIx+TA5Z6yg
/Tzp9Cy61t/GA95mPOS2NPRQ/RLn9T37QiwibdXGEWFyrEVLDyRO+RKV182IPQYwpgQ50fTd7Z4F
9yLNafHtkT0iBf1/O9vOzKQXh1FaeDY/8sNXHttToXRxROmdU0osBd8MqTALxZQ6+GsMuKYGcFxS
v2Ov57kaLfuJxdg0KYQXl3v/oPlAn/m51Jxjdjv5JFaFSTbou+CWnajs/DKcJbMP1a41wbqyxj1a
jx3JqUDW9EaKEHExqcbcDxxR4uwPn0f1hyfKjQmLf7YwVKJahoFxAhKTu6fBxt5HiLLZPX6Fj5Mo
RbFkDdaxaQiH6ARMAh5/bCyDFro1OUs3ZM3Ap8H5KMZcRU4moI3mcWcolumShPfHEYai1somKToA
kBtR69Ymp1slSVpXMUpKRwYN1R99lmfgTyoXd4vJCHekcZ6D+9UAmTMTV+3NrkZ7MtwirIHikX5l
TTWtzqV/nJZmrBFO30/zzAoRwokOiqD0iJp0Dg1wAPT/WiaP8YIbMWQGYXeWkHTvVqmIO5cAFmPc
kWs+ThaQ8jI2XpaK8T+va7rMgOD5uIBCqWXP5pqH/GP7BMGbl+ibn6Qu778UszvR3rcMiliS0X9R
dNegY5Hj2WeWWTkXo20bbvZ6fX/1tpdhRAJ+xXBz9wcwriatPP0mekzq6CL4UcHKFA5Wud5qityZ
ZtVg+oNzfxvvCdMAUprodETwO7uW8mDr0G/U3eWvlo7AIn1WmLvfHhbQmL9SfXFEDpk4XLdPgAqR
q+/9TDyA5dyKdZM8+Oef7BrAlyyHLxSAwYDQWotTqGk9cSYvORAcwgfPlqPMuxvXAUycabhSh4ds
mxb5b+ZLzQ3QJSMeAmhZXtMfyZZRRDKJFGX26VeeeKMjCfnj3xD5uWzMIjW7LS0DaXSwwf0owT7V
tKe96zfD9UI52l9v+25ETepd/8nObHzsCxEiwl1STyKyAiInjzHNlYWLM+8vM5wf1lqN3W0+ZEvv
GWFKTJCAc5c0UmUGt0lex6XlGFd3yKZvKDj+H1DHJ4/8kHO4XsYBvX+QHFsgBq7vnIe6MKZXm4Wo
1HFJvUa2Yo/HKU6x71mNhMewYLov3EjSlJiHIwviQWmiJY+16QzzwNNjhgVtiWnnS0lr0Zy6XZ2h
YyhoJrPfkqcfXta8BqiBg7O5HXGH2MdnO1LNee9PuJtxQh1BuxOQfNX8u72Na1ykGAxkW4HOpCl+
mOxav6EzW0rMO0mVgjeTMUQc0lDuwbcgdaXflcto4jit50tZQqaGQMH0Yz8+bFklplqnhl0vVmLY
9aqZFWDvm0TFJkNwR1dSh0NTzfEk/6bLQke5y1NzUBYztxLUwJrNupBZ2fZVXi1LY0k67IlxQPMX
4NgjaGr3saqYaxrI8aoGGpVyOFkdfCJP5flB7KY0fSxJZN3PZ6mZPHVPnfBC3xIDalqRXxeDvqWk
er0RybeYRSkVDsMMFE8FmP6ka8QzghT3IO/PdWfVWxXBRIcjqa4tG6YEKB7nqqqCY1nAyo74pstl
H3NsSq7bwvfgNXluoaqEZzhAt6NxWtGMFDuu9KuqPAvB2rMkZtbxsY948xKBsXn6SYteB7vEHH/j
I8rFdX59F9n/pnRmEmkNSV6jCnLCpPFokq3seHObK0djrDmDuRzlzOaxSV5Wmeyg+y9tDHcKs98d
+6oSPdy1ZXKYX6Im4Pi6gZ7CyN+lPA5okJx5JanuGR+s++qS51Vc07wbiXDZTea4Pg/SgCBEpmot
TLuGDehHMQBN76EaoUoIT3xVnGLvlkqSP3nUXM9oaIMBfh7mMBSJ1nb9YhTdu8pYAYnFiH2Vo/6Q
ADBLh6Knzc6g+EPW5UJAtdSCQmbsNn+euJtShxSzRa7D72xsCpoPRExdioHngvHKxRAhdf8uxUb/
UZfGoGE16NcKuAJNbCgvi8d/bwlneMOOp4vmVi5huUkUDepC8J56fEVZn7Wi5sX0amGcxuJgICCm
mx1kml4DL3SrTesiLxtl/7pkpymwPNPQofFuppu13/MWlgCp6QGLQnMys8hbnnAGhzZPG03hmxNG
N9DmazwNpPJkmJlz8TZtli+LLyS/rWLg5aMe2DSlxstdso3HZ2dKok59PvCDelIE1CNuhgeUBmcC
dQyL+p7J/s1MYwB3UGchyQCEkQHdSwwUoLoEDqHXvkQ9FXkfiT0b+A2D0xDEnbysT0VFmmyBCXuw
rBpLVzQM3QbPs74aaLuK4R9F6FrjcGR7tHPCXQa+UgbAJs/3Wsomm0kRjrVPVD1I1G7jj7f/uGfp
A0Cq0wOqwACurnF7cpAcGR1QF06gVni3IkoghjqGgUH2y/hHraTGkCjODF2SrRYe1ZzKW1EXnPSc
68DymibzX8TooiuueTSUhxDfYJMnIfPwTBigJ0b9rVPF5MFpJShLWdzp5UP9js1Qzn/sUJEvSODh
CKjwsVM61T7WAprMG5SaEL2AYg1MmM//wJCTaUSrwa6KO0XzISCmkFoqIiZorPn7SY0ej/B27pz/
wfQkdxDswm1WODOby3yae+Z8138n+Zu0nCEmS4mjy2O6VXZHKnaxYWQgVEqL4HWRLMAQMfyZtNfn
31GeZSpJN3xvVV8uqDZnLEA5xvMnOwfeSkv0H2GTnRBvZz6kIdyG/YuA0eowkAkr9VHR5AqW20kR
V9BlqZyFuhWWpleeeenIVs9KnwqMrK91HyV+l+HIq0Ob+v3FgOIahfU1JVz+g80nsZe5OK6L4Es+
9eDvsLlJS9Vua8SRDE+9Tldr/ejWx3QVWmiyxMYA2IqoEtcUMK0J/hDaEc+qioiDNg0COqW5CwMv
Hbo6tIt/W0TIJFiLp6iGYSqifefgvhJz7CvxWdM+o9TIbWP4QoBDl6s4RauZqV+T6AcXONXr5XQ0
2D7sixlK0u2zgOX8gg9NzhrjLZHNiqIiMWZklK7TAYOyH/DwT7jNeT7UHRdnAT4d95Vh8/JdGDzZ
/PlbZNWZR3i1TwsKqdNBFGlTwd/523DKNA3mlhUE8TkqgJFTzEecm7VXkejV6qmPhvtdReEY0yww
fucJL4vsxsIrrhmh/VUZukTpMmUXeMkW1/2OWnTgd/1cNOlLz9xYk0fGysYUYToQn/8dt5ke2MUW
PfkN+mYKhmZnJE8pP7DlleKVlwj9W0jQwE5dHMCNISKCUGhITAcSTFyEHZ/GL3IVhY2vrjHpKa2U
sNa1Ye+vWuxVuvcoy4nFk8kbYX46ujuxonEg0ekN6u4M8ZJ1uirH11IVlPSoSykDSUeld5UvdToO
PihU6cg1pcNMEmp1xwfDb0dhkRiKoFAXPdCc2V3KRMa8622ctBAE8zTEJwIZIyTOIvl4vbd4MmYt
SyrFLaMRll5un7OGWKNPdkrCigrWL3dbRsfFoHj0dgpBChc3QBi7J2W6qWaGRUP6E4ejLBn/qQNj
4Ql/AF1Swwwh5nWlrGFhToQnKaPtPZsOPfhwJo3oM1RkWXAqVf0IFssunXmF+02L+bkPY4rfCl7R
ybdF66fiT16IhoZX9068hbz0AYCBJr3kOzAC8RHuhschJQ3qDmJirxk5rFDvs+VsSV2xji4qEzGp
AZuE0ZidS4yNXJfvxfAGPUAMRQEegJc7q4IFmxhifVF1lLXhB7XDUmc3IuF7s5wBvjWnrhdgSPn3
ZQJCqEApmsTwFeI8lPY2SbEC/po7LkALuAM7WFybSR4mwH1hwFQpLRU3Z/ZtuaJ7wYhTJ9m27UAH
Gu3zXc2r6O3Xcn+6lnzy11ygtUiYhdUvzaQvEZKR8778Rn8ICMjq3F+LINIJNHYjDjUhYy1ZNT+7
VYa7hHZCuP3qFN77V9LJ2yXzp3J/5fm4lS1gb2Ol/MfKRtqGGzpr/FP53BX19TgLwr8z1XYqoGtv
qgXtL4UUCdIHPgdvl9cOSRzQTQGxHa4v5HyYgM6oj6AUcYups9qAckQzlJXqPrp6DazeOGtW5BQg
cPWbJ6safbxmxkp3IusUWIdQgSrR4MiJlLiTmfMkYs3t3qZEJhcQcGEM8+HMYHy7F5105Rr9FSZQ
u2Idm/bQAfNansZLaWcGq7Oj0wA5baeIp7endU6to098uht5m/BRKoDtQ9UiaTSoMCv67YuttnGJ
OHuixwmWm1ilMsNwZk1xIF0/29dcVQSWl4UhsM+e3MVZbltfPLCdMsRSkK+FmLQPr5xhXHzLXK81
iyxic/A8ps3XZaKFV+dwpGzGmpq7IYrkP97FmS/aRD6jSrB90A5NwR7ZhnH5chIvWVaYlVH+r70Y
tTP9ESzAy4qZREn9jLRarXbV4jcrPZRxmMiyISFz357v/u4fzSNwozEXF7bFDYe4YHriPbKQ/ME/
Xf+wdYlAUeKeA1yNkwZoAqFrdeuQD2HkS/qQiN2u3/YTjRiXgYOCiaFUJM4R5a5kOym1duySIdU8
GOn99o49ySZnTRwOZcwmUmAwkfJbJ5PqnChRGKOjg32asr3mqsIsU5tmETYYHpXsl0p2uVJPMlSN
qPTVreRUyts6+85NsoMwiiNB1ideYeU+/CJxv8UZDenivVra2+MziJUCcwnFxpiE4J61DPr9gKFg
qlfnL8/AwEyIz2/ghjKHaVhrnLOFvlOq6N1nTypeaUDj08Qb0ftl2LJGIUK7HH2/ixT8++VlpIoD
ZNN5xDxyi7qpBoIOAy3bQRBUsoAtGjdKfaGVHq4O2umoRPAZqgOcJex0xvPg9A9I3WRkXrk4Rzmi
tOL6YsPsxZZ7OjKc/5Yt/XmihetsbMpNcXD4Vg3mn5ht9KA1ERYAykP2Fin+2tH2JmLElyyd7IqE
tZWa/jLdxE+PG5s08+3hhuCJcoeaKF6UFWhNGJUbl8lAQ5ju4DxaNiihsM4ypXzxzir3r0oEmTKy
gTVRQavL/dJ5HBDbKy1+0xJoIx/EPNkChvlwSMIVokWivNgz2paxCKfm138yaqbDKipOHiO7nkJn
QSIpMOWauwdtvC1R+aEbA0juQ6dGlQhAQtChrl3PUW9OI3EYZXNjM6wZ/PMC5NYZhLWRTAow5rGz
Cd/5mLszc6m2kH7tjN+7HkSeQD9DeEjjl69MqO2W+N3CdcE6RMvELcjoY0JnGIBchfnhd8pNl/k6
G9hEFJAMRPqZkynE6roPh1qWVhOYpwtLT55+iZhZMN8YtOUXb+X0dHUDAaUuIOdkdsvH4RF4P1AD
G7Y3hS1tmw1XKcRgoHA1JU+KP7tWbLpoeSAm2eXDjD0Uokc/lGcuFvCeHfunpNWpeSPqjaIQoVfH
t2iCh/UgqKI4pjbVDlfkcZp6jlTD8o4ZrpGGsSCWsvJTd9SXNzsrmvaoEl/SbpzeSLKRXgypud+1
bzaZoV3miHhvxzN+Mel9NXyRMOiDPwQrgx5Wo5G3U3aYNGg2RQInZocMkVBy2Il6fUrPLYdaHUz8
FvkHxOj0ZjCx6D56YTFPm6+NvBy7uHCcN0VLamOUD19eEKXwM8w5+nBX+bMSYNlhSspxBFSEAovn
lCdx8OaRpSzEYHAQS7hq1wLW73D93361Rph9EsMoKtdvCVAHC+aghSPbjKoUw1VUFOJSTCokjx9g
6b5vL/5tJAgmDGq3GZDHjCsooKRIC46vJ47/cjRx8kE13MCKE1zhaMq8W7ZfEnUSu7kRECAbIVox
PJbKG1F3kkVwztpOYI7SNSWNeNBfOyzmRPgzFa55mQiVBPfzjaBmNMQ8VA414cZITMypo1mFPRqu
hQjOmOmaffAXGrDl6rb0cq7kRCaLfu5aN17+zk3oGcM6Wo6g5ccxhZACs8GQV3RLS28IgQQurSzT
MV5sroCUES2RvpNTg3pjMWfYTgCckGUKAw4RMLXrra2POduTN4Ci2g2wtuIAhk31sQZtfhmu+cIO
wpqraOOhF7Xuutr62esMN1EpMo2SHjMJunIwnUWLFynAs3oN1jU8j+ez3ADJShbiyI5VKJCEHbXP
D5RbO6tJZ+eNeP74NaQEeIHjRUX+Lnjee62pdNUIG66gNumy3b/qzHPoz4Ea/oiPJW+uvWiFAA46
nWnl5rhA+NBYEfHQD1vzRGhV1JqVEJ/gx5OTlyos5nMJG4Pr13hJTQMkFbkONPvBI9k1SbYZZkiX
C+W5p55CW/WmlBOX0CIUrSNFoa8bTFBxnlIsy/4WuG/4koDNs63p1jBKoWow1Sci4iHbyuseCSV+
Ls31hr6BydBbyhA9nTkz0Q/grb2r1tZGfo/B/Gtk4jKzRI9eJlaYHEtycTu7okf95Fc0sqDWiLyW
7/iEiiSnWJmAkALIxc/U2zCbpF4+C32nTT+ps/C3Y+UkcI+ZK4tN/NtmjkU83DC4m3uujTcd9Li1
jk2VuCsoOpOkuEzTuaczJMj0WZZd3d9zH9u6DNZHlDEZGc70sjiXXz8QHqsh7zpDQSUNxuuD9sPY
P1KZxaEhGei4kYWP5zZAZ8cCf3gntA5bal5618LdNiggF8o2EOtb7yHQpt2fV4r1pcEzhuIkHQX/
rs7T30FuElKtO+23lt8qRIynTuqIRCNc4O56mA0K4PksmkXP9YwSmpkq5yDUYrC2JHHZlMg7hzvw
St8Qmv/hEUoixFXRn0Vx9kVM7m01sGoxYSu5bgN8O+knsmsbJybQowJjbQQpcYWK7BY4jJISawSd
w0wXd9nyfq7Ygi1/3utK4IA4xXmn7Jl7hsi3bk3Z+ZzIR1edjgZAVA9gYPTHXd/lDvMUgNmK+XfU
KbY3PK0e7pB4C8dNHY6gNemCZtpuZbEXMRbgokRNpXb+NssYAlujvVWUfb5Dh3RyTVQkCC+Y8QAh
jBS51G6Mbvf8bBega1WqqngkMYBZVOL9HArgyYdJ0meSqYoy1R7xE3Dx3g2WM890wElmphUuL7+c
8x4TTJyVf/iLwBojJY42kZKaIgv4eKyOWNoVLiEiuylCW1DWlKAf7CrMScryWGPer/B0f9PEpM/I
rt2G+oKQyrS9INs/3gzbizccJyBt6tG4yYSsTo1Hq7IRj1YcMdqM1fkGgEFiF3INa+ZHak4ofwsM
jxuCjVkreAdHb7nedoB0pmjaA61BNwKbv9AHZ15Ud4KXLtbxNE1qw7lpWI/CdABWq4gQSqNFo8jL
XixJqafGZqgs8fntjkSbjJK+gbS0dgD6VJoJGmvAc5txehfl6o1m08YDR6sc854lVzEPwy9yrVf8
FydlRyQsQ3lQ+IcqznAXBkgNBl/2DwVO0n6AAoPC7RbIQdqvboYqliKJEQTOB6BQ9tVPoKofSS3U
v6BVDgSCEUdEyFM5YKAekw9L++HDvLIsExLx8XnNlCP5I6sFU3IRzF0XvGFYatUJ0rXoPpiS0gK6
j0IpSoIp8cicvJB5H5N7y5NegzvXZMf7mY3raCrKEisNroeOEaPqaD+E1VzKlBThmVcQYN6aQUrD
CxaHA9yT629JAlQz8wjetWisSQiN4k0/RSpibI4ugXzNnjbvQOYLAcUWW5i54WWBofZh1PFVVKk7
wlLMp9ljb2TRBTK/nDuPVWlz8pLYpUGOhGjU4uCH8uF218nUnQOmTGy8QDFWJ1Pi5wkbmyPaPeB5
riLkvwUco7wuGFXF4sh0f+6AII/FvDuP8T4xa+1qoa0cDRlRhumKf2tqlNccE6X66A2+yYjP9CSk
Hveev2VWxsOCUZ4IwBD3pv/C917RYfeheCwf3LPDKzGdh52SLvpsuXh42LFbkpF6nBwMBFfL1GID
R9TNEcA7fkpEV9+r6nK89Z3/FlKehK2wVR7Trs+8zGcdWEvlc4Px44+lLu8s3sRQWo52BNM2+J4a
DTX+gT8A6ditG6HNkTzV0JLnlW9GE5QLcMk0GFGk5WIhHogyRo5NSEjpkBzOM7QF/aPAQszQcG/g
j05ycY+zB7qMDtFmFOKglXnf/3z+Ul7CQyWe25d75dSbQcrgxwPDBQyPtsT4/lBtsVolKR9mBsq0
uRkoYlbY/aRqGsdTeV4WOSzDM1X8BOmLc05ZXDEzvi7kiUQKWZ1rEvvNlErZSejdG48CBeptWMXP
vBu0C7clAWa/0VCL2kQ8dUM2tXF1h5PkcyUw9/WSPnL487GZ/ZRU8QSIgZ0bh+uhrW+FNXZ3f6Rj
6jYOu0zk5kYxjwAzuixQ+KaYk8whg5kXpEIytH4zkjtEtna6m5fUpio2vINNBwBv8Zt3X9iznWs/
ZGeuQ4bJFxQoly/CgtE9FWtkrflqKTtu2r6OZZsZzOSFA7d+NiLGjoH2JxHsLSEjR+HIevdB1V5z
m/MHeLWGMrkjWqvAifeJrm5+YncYPBAngNHLbX0MrgCnbsmMYfbUgmO6x3PUleQSx7jiZkiQ1IuJ
tjnBXVgn+uVVKCa8hiFhY7C7d4k/TAYAcwXh4UmlqUen/NpZ9Up+bKsszpllImAGYPFFBalnHFLe
Apg7n5zLfslwWdbPKPRf8BfFIttIA2XuhKXOq1XI0j7K43+HH2SQqtoqc/GyMXh2RAk5DdnJKz0g
ZIbKqS3eZoCR5RDNr9ZbYjXiLkegUkWEp3yzCfd0nFI5EkgOjjC5FjO4R6MJicb3SZTCxUpyQBCU
09GFHCogAavPt2zELifAXK1cTkkORKC56zd9RNRkSH8IiMLqam6Egwu2z2R1HGWPbj0AYdzBvZmN
zmPI/s+enO9mJvW2RmlyAMnV3HEBnqRwJhUIdeVNe+UJ14k8Euvr7gSoRSIKhx+xyVyIaHDWTwM+
YrYFqqHYlbZkeGP862F7J9qZBJtgsZjgmuyq8fJPSrYvbfQKeqTQ0gHMnzlCPpErC3Ak/nYV8JYb
4stvZQa4yQVZKtiIpPtEjnKsSi5dhDbVPS47FqpvEse24L5x2kBqqK5ntg0gqYnXPTHq62pWXxYp
t7EAk4sAamgtkPBzyeRXW+0KQwTh5JLk+8ocYhYkfJX01kXSYuxNCb3K3Nq5H3zoGvww68XRIfsW
JJmtUZE9a0Gl/1izH175TqNbWYDgzVta+fhjvkk1eQHHSuZsBUXFaVw6ynIkl1z2Xz+bFNsN9dcu
xpsQ/fjsJM9280QCL9dZTAjRxFi/CzaDAshZxUFGBMSmyfOSCtgZJnUvHCOxUpBDmDmp8BUsW2rB
b/oxvKzKXAJD/6WJPwrB1E+T0F4JmC8MgqDua20aWAwSsrmFCt0+pjHsGDjefrbhRhvNamSxM798
HphUiwAwe7QAVsiDZb3nM1iTdpkXQtMTfhfhxw930u1kbhtLznwsvpROMqzY55H5eDcGUH1c0IDl
zAkufck9nzkxFd1wMKeNwBg7CJiFFBR1ieuWZJvLClN3Hos+OJeKDtGiL1P/+5PaFqrI3lX0J8rs
QffMDX9nLrqPk6D1u2hL1cpWYdsH88OGq8Mmq4MbRejVIRZCO4PXzG9m/KxoWlvqUZzuDV7GlJTa
fKFlmuCJymsZvDpvb9N6jROOxMVd+W1SSlBG3MHFIfVyhJyMwsY2X2Psew4/OrxD3BNYrGeH6iQL
tMv5hCuS+ad0SrqhyXQW4TYkDN9RUlc3DoNGv6U2sjrC5iXBLtULFl4JibOEC3bHUSHXgD1RU3Ru
2jcfdqv4BnFOFWz8AJp3zVvs3MHqAbfl6BcdtgnIIhTBZ0JcArxf9nPj8ug9alXXA58U9nWWiVBV
CIzyLuVXSPz40fnlkS/svlYzpStyGXAEh4uJ5UwnN/Jjf9ebjyHYU0D0Ahzs09ZYpoq1tn3QL4V5
/xOUOJIuk9wLGYBDO6y7GOI26TG01MEUWfyjaILz4OW9LrbaNCovhhVxatUJxbO+tOq/fn3XnfhA
S/MTo71GlNzrjBQUOZj62ws8+QYnNnLorK7zzDyf/BT5Mivj1p4J1OG0a5u3FVjVa1GLU0o/s/NX
cCLvD6IJw7HWuUeH7A5oQKk0zN+xrhRZBswGn41Je4DWX3AEOpzDEVGuSINPdPxe1zTdU+HhGYH2
7SNT+/mF91JEokJ4alwGiY9LtrVUPgTpZDq3ENTsswSLUineM8JxE4jvhiwTPfIf3DFuEd8Y3bvo
kl5AtFhjp8h29mWVptqn7dzUcvp/s7MAgx4RJWl8eOnOclKrP4Pv4Ee1BWkzg+q7xhCDgxBvdXM/
bLQslsjL/s+Zujw8F0TBfetCXwWf3kVEw9oy7y/dVXtBo3Mlk1gEj8IVzzJZ8oyMKjTzRrVuWTx+
07Y5MPWtkykcVrVHwwYcxMRAklZ5IDcIaJenDTwkek9JeX1igI7wTIkxTKxS2tqzwqo6R1PvTu12
XvZN8pzJt3EoG5FgyPV/i/cFAUB6A4N+29CVFUEU73BAKg5m9EerTqPZ/cUd3WC1XpPVOND4wj+g
Lj4rRBnXeIchKZh24lUGBAmhbPxhqOE0kJRXKsyAJjMUe5fi5ptawW9J+sWLIRor8uMOuHFmTU+0
SZAALpalaHW/G7ZZMFDj1N9deDxLel6Ye6gobZZpuo48rv2hCeYPlBJ1l7fk2rvYecQO2jGpa3Hd
DHaIP2PyBy7mju8q3FUMh8E1hXgvVNAd5UirHknkFroSEByFSiHbmlhYmhl5WqB+r3tz06FZ8UeS
1QPJ0P0wbg4JTdHbox05sRlAn0uCQlOSOLLt7cGtm680iZXy1c6Exl6PIMl/hQYr0jnKImjOfabU
syW9SrQuV33pyNgK0HjKW94LJn2ek7RGCl+wB6SDNQTxM61LwwSQRXaamhCMgN2a79BIoCZCFVJ8
CnXBYxMgluDzP7tbFIEu776uxpxLOAC6Ta4aJipWTFEZpdpONWe/vlolAkGR9a0XeMNhMioSye+p
Nbc+nQbaE1M5m7p14UGLtPOFzv3IGlwCdA5QB9FJJNZhrMhjm+mRuJbxQBTQ7BNSgaDYvaH0i4x4
doGI/k2wuzhm90SGV+P9wIX0TBevuomem8xs/H9K5oHgPX//vHi7MqhbdT5a0jCiliPtDdKKuNPo
tz/YCfjmZvMMnsEHILG4IgK4wLcKSlUtJRbRziQMuifrPJ1ipkANnbrdzZVBA5B6KKYjObomhfpF
akfqG3wu2yR2s+yYA47KCWTzd3lhW8RsZCLokEepYiCMWcGJCPnd1QqU5Xgdu62MxGF2+3MGBOuf
afzVp/B2HMSneu2IS843/IxL8Kt52FzzTB5iX0sWyGD94nV999iSw+9E/u92U+Jabb4RHFo9eyou
IJNohAay1tDU8Jz1HemNxhxpLLAJCOvHXJpbGQ7DCWS556jb+x44TzV1sOCZ5i1JpEn9X9bUpqh+
GaAc1AyAqOm9ouQ1d3WGLZc++C1/NkfskYDEltExBgxk1t7+sRf2eEB9qOot0XtYIMVwcK0NFQrD
UgVBnaiLANk23b549zwrDy/fJmsLU4DnAILfgIDPORuOMSjt9wtC0MBRAwUgfmNbrbgiSQn75wB3
e9gNszezgEdkRYRdZJ1iJ/tFICtrLC3Gf7hgn/VhiWnn3P9/H8FMDSuQhIlHMwM6afOvxPT18vOX
ve84DCOOF2NmPljEGsK8qtmCkEWCXleqC0YdNuMedE6QqtnHfIMm9qRxU6TKZdSolFS3x8ncyN4J
0tZoSx/v1iU3TS0XACzm+LO7mhLqchwPm3fYulD4MtjsPSlkDuQJDoN/N2DIJNHfUnZAEBDHv2YR
tI97xCwxUpf+aEpa+Zj9G2lnfseV+XIWbq1n47vPqd4rgExiJ+vhM/gyvM1GhIFgZZSWG0fmp5p6
nJc9Xlti2Fc8JWYCPf+CD41dqcvqpGPAUUXFqtd8qmgnXpZ6TKkiQ5CI45ywB4jRhuBsuuhfwnVe
h/eEkCExr+hQ/ryRLqaaEi5ADHGPtlGovV6XEjCyEFGLgQFM1I88e+W1gkNk7VugDXvNZOI5ecQ1
Uy6GuEKo9Miyiyso+1bBh9ZyZVo3SKxqDb/uhaYBHHKM55zIokwQ2sA1DDJec5/Sh/M/DnMOE7J+
qaKeZLhLA+tXcODtgGQBVixZ45MEay8n06lWacgx8qYiZ+VuKm7lZ2wSr111tnHQE+yonufl5J/W
c3wAC3wG31PT7ukNWX7NTXn9PNcUZ3/NS6CVwbXyzeEUsS3Wqf/nHoC5vIdUo48SqUa/1fsaCF3o
DPDJqg0UrdjEtcw/ZWzgoFmQhkX3OExd0zdQSmEUpro2XDp25zY+NojfHUHVRCo1NN8iauCZSc+q
FO9eKgCHoRkuSDNduDVNs19M5VoLDFr+FBVayqoc8wPzKi+Z4WVWX8WGa6cUhBXhR+q7E2HG2mW0
L+tYGscIJ/k5kT+aM9Cl2e2Ph3HYHahdTUR06FinUNekXOtTZpg5/v8c7PB50X+n3l9XTPDL/pSH
JTnhdtEc7QmsfRz3PxghyHbJ8LdNMVsqzh7PIRm5gdwyV39999c/hLdxBhnBNoJ0bbjwEw837a82
LG96ER41hVMhJBfb3Yy5PNOq0cmKB/TcUlbfUZrZbC7JfCugN2R7JaoaxcSe3hw0F5MlGOiP2KCx
nby2HqeIHOmwYvj3m+SzCdAOHDWxrcC54K5mWFUoIwDX6l1rEbIgoZQftwUs+Wjd0H9nrLIJCSWi
GuOFpHGRlXeUVJevMcC2XWVJVTldwSN7YZLbHEL55fDpf2jAW3Lz6zpCYIWUcYyGmgLExwNBcFjb
QxgaN4Pz1JFjNo24LlXwYoxd83kafn6o2MI+8lBPt+lEiYPdipD7vJqw4WYK9hOw3u3w2g3mVUgm
NKkQLk1PHzS6jauJF2f62LRdarwjb5iCUXuh0yQLpxQY6H9mUYhjgyDwZ41EXk/A4tFFLZs4JVD7
Jw1zujFozV83LaxhpZhw8sZlRMTC22doZljKyi6USU4fjIQNfi4v36l0XyiTOmDnU3ogLmKVtWBv
KOzrJppogrtdZOYzBC3fKLP3+Qn8+Op3Y/M71fqUj5xsSz2ykaYUnmSDWdpArHUN54ADbGcT31FK
bAdlms04+kX5lyaAl9K5QvwwVdK13mE8di7trkuskkOBR85rRVIckJNacmaNFgUau7i5td1fzDeH
7/u1fk9bo44KCs831RuGeWEoyYfrsX5zra1jDK0IXw24WXKEYXIbpu+LZGgGhDylLbCUjCJl3rVN
R9RqyXqWL0iKIqC5P8nOL84nQ9Q1naTpr6PJqI35XnZZl5AyAH/oX5a2nbSIY1uF7wM4vS/wZr+Y
2e27hiIv7Ttisu6COm2Mc+k//4RNf4Y3iuPhi6atqxfdTrCkxfJcqYmL8+Zq+PPjzQTONyipoNuN
kquRiqMtnTxX8PoIBftxAVY+uKsJKqG8Rwv2bJ+Ham8KUbu25ws/fh61DUHNqFUb9O5x8VvC+YGU
2M0fONmb73h21PP3QDZUJiNUSvh3EN+ZnvjdS9ijcVzavF5XK9LVAUfgKuaRIdALMfaWC0FnTaRO
F+N9Afg2iZ2N3RD0KWhsI3l3pDo4dbxW+Q7IJfQMe2ImtLnNJHNBY3wvybTa+z4dm7lkRonptgSq
BmrAF1ItK0hwDJ3OxxLeWnvMtQTUmLr0tK1fo0Pd6ZeHqk4GGyJz0ZNlTc1zG77oWE8knBagBBkJ
LSqVDVpo3t/5KIKhI/aln5arpYPm5kzoJNrWTRbyUxZxvoDyF3x+7lRaeSM62qThoPtm29KFzuXi
0BVjB5CsxSZldC9HvMXtAGbImeSW5hnQEy6yKIPqmCzhi9MNl2DhU/RTReJH2nv2EWQ6sy4xia0z
bebJkqnwZAezVAVHcqJwY0BC39jvuQpKexgADwQMp7jKHnH6WxKyh2o4sD+pGu0NN21HlOshYdKR
kCYql0uCga3Cml89RKX2vviqFw9/zikumQ7H/GRBv42IkvYt/Qa8GIDTtYeh5IVnDgx+XLmwPSx1
olRKFJ1qT7UEyZfQnDRZNDBkvGxy+M0i517uaurmueqdCltJEEBE4LmKhlSzjYiJGGwOc0fdiMK/
F6SbG65dHRFUHGt+/Mij6lHdkbRbwv6KQF6WGpljo7JL8X/E641Avor5cAydEZ+gkokG9w/im568
76j6t24zFMiGK6RjPg0Dl68TMsKthk9QOukPXs7oi75pUhjL6qZG0uPb+zyffA2nZws94JsTT+En
unq+ErBwB4DXtyfUSo/1b7NCGw/VnVPczZgQYWYDP+fdvm2Kdkdl3f/T310eKSDMoJggo97MDD0f
GspuIFHYwKYf6k0UVmvtVZypZJzg9Pi48dyRQs89b2tqir1rIzAz/ZpMX/Oe/4jzKde464HwQBDb
Xp4x41tQcftdnYPnhNMRyS2HhJ0xSV3H3SEX/2D/zixnmPU62gYltOJImO4oXK5rIin7O0Disb90
dyJXBJVf1RNy2TUjOykVIW08tPiP8UBFzygx7LFUP37tBZR1dE8K34YqK+8blfGBrgvn9CZhyMa0
caOCqePc7PxOZ4htqAhVHNiW7EqrSIFa06O3r1edrkyvYthsbcHzfQDP4x06XDwpVWN7vVHUeegZ
AYcsyKWs+KjQRQuw1OjKR78ZTYqyFPbt2wyTha6z4yYKXt7QbTXj6vReffu4WuQwNkdSxlwn/rI0
iUDegR291i9rWOksRMjH03ZSdtAbo7X1rX0b1Knzoo6VlpO2wuzREupc29PEnopl4fvEUb+Io4y4
luoTlD5by1uLp//IWPMsAUDy5Y3xKajgQjr9rJtjf+dlUmSqb/eXUcqd7+rBAvI32ueTUNFwrSjr
hjeGwCjiAMpMCOrwJv2AfgOHeEO1QdlgiVfMxM7qhwUXx0ES/wxfOMnRGNmBha01ohJKIDooruqV
TBMolmoK0uHMvVHteupgvTR6vRQevyD3U54Eb3eI6+gWNqyds90ZHdMn/qwv/BXS2rf4dbHnGVHL
FUnsJCxiThnmKX1fGdiQVNZb5TbGfubcQUuBE2IbYERyctIKCuv7JfhXHeyVycwfJgRLHO/B/e2v
kFsRDdzyxYcqwGBeqA5Td7tTjRCPB46D42ag/+M7YvsS8LOV5yM9CR2kf39qKxtXzTTb9geH+nzI
RlmPwPwLHgTjkHL+sjueci7WmDSYo7ZOpyi4BW8F13lyMvDbPuRK/O3aRiTUTKIpRg521vrVrDB0
ssayXH9BXuCB4PC1qDqYJJ8NtUuzAylSwkxxuH0y2h0kBIcBgRcPztMBncojv+y9PaOltT7x/EpB
kTDDVk/CMTX4NOmzocQgY/q8j5cp7tMR6UeG3y01M0aizfUy7TwW5JPxiSxzJTtq5Mvm+lbXS4aa
3aycKuwkHW/+WZQ17v9k/qaVC+UVgsVRRRbEj65rdkmoIrPeY62foc/tjWyqMe8k5KjY1TzwUInc
oHJPrIzPsFj9NJj0bnqeFw8JY+zb0mEVGmfSLm3NrehJzAmuIZ62ajJpi9Pg7Og2DjVqKlS5LXmv
2xi+A7Nkps8Aq805NKGZBjro3vddd9nhxRX9MluOqDLtQLI+0/WtEuA5AopLjrC0jL42oBqeVajQ
nQYEMSFkMkfOiS2V/XIiNjrCY2lyOljthZ4Et7ZHVOz0rg6CIa+McybS7WCKTBq3mXuURZHD+ypN
BoU2uLU1J7Chg3YWBqa8WqgB31Qy6P4Gq/IXgn/gd7rZOVOmlpTE+2wPMdhL1OX2Sz8jOsddph5g
i+sExyYZyQC0GhHQU86wEMT7cd0bSfgGXDb+7ETBNBEVAprV+gDNs5eET7JG4DABpymw35XTy7wb
3i0mCTGloFPFqUTJJ+e6hU/tFYqDBATirpkecf4HrXCtnyLvdfqQvfYHjKMi9pZVhrO+fUBW+x3s
8FN0EpgoNK7qrEpZmGUb3TcnINsWdeMaDe0MObNT6kyyw+EklaeFXkZCYnJIrJ/8vpwPJMObDxUw
q4GKpN06KlFjmwa3Ab+RFNJa68YJadvlRiA+IXlppUOGc1mZk3QTpTJs3EUxoio2obmO6mrxJ1Mi
rPEhOZCO2fMyNe89klJuuQP+APdUbfwuQz/0O9fcZcEvGnGZmgNYhnRig5z/YdJntEVgNrQVor+M
0gB7b9HKUdnJ33tuzBVGu0PXHZLJ9ZsKgVGJ1ovZ9qjvQVz2amR49JVu2Z/2zJVroG6f/Y4Fti6o
dsxLP82M5ZDgFtCq0u5uborfwsukQlFGk7H2oiR2JIUFjEwdvMCSFnnxPblK+VWBE5Gx5oF2Btd1
3rIie2/OKQw/m0oxhfKNXVpphe/BUtFDcuVYL13kbHja8xOJfNtuVGFH/idw1XSy4U1gPvauNa53
I/ViaU0L9BCffclPraGVOVugruT48Ipg0EL0iLfpXUIrDh2pN+zQxbwZW8ETwqOa+8bJU6QBzMNh
OohkNRosc51Av8QsUylv3qECfJRpwpeXYG6iXLBgSXKEtUEg+Tw6925Uc1E8WxKreKWzxw+DUaux
d/p83x52g0l9rcHltOe2YJxMJIn+dBAYSEjlyvWG3DXyvFQJciW54FBPw9D14xyTlO2FfpQnU334
V3ZQ4X0KR75mySCKFXmoRjJqrLXCrBWPHWQOS2NyRvXbp42uShPz06HNJqZ9YUphUncgWiWlqS6w
JSqXMQ3vCeSURMhlUEyNsGKXc5/8IMRlkS7rO2otmmj72Oc+Cs/gDlxG8YLjgEtcyIzm8sLbWTUX
FSqkCeFz5TKOol6PnnBqeAioZ78893sNvNCLbGlzVfYR/p32mHx9xjaQhtTlY91l6ekZ/Y5MsQV2
P5nPE8KorhXuBN73t0lFA39glavy9JdaF6b/apGiiG8kPWXXSbtry1lM+uGKrFXrc0I+iENXzEAo
/LZsNrPBwFGoBjdGekwwa/IkabRohcI24roP5Iv7IYhaIyeWvpmeFR7OPoQNY3mK6L1dIhBBH6ub
E3cbn6zLzlEZjZuRzLNRqTqMkLKTM3Z6GvrcUlsNUk9bHG8/RhWJofsv75m1nORpIE/zDtxGG8IL
lb6LY84w7sFCIwZAWOaF7GXxLEnN/YiuTKzYsu+8t1uD94N89QczDZVtcorGytdBUAexkoq1ZhlO
vPAmgJani3x9BlWevLFUT7CMxaRCCANLStM2es6aRkOf+6ETS3whJOEwesic2M444phLaW59LyQ/
si92Qny3CrIrdF4VwwUVkm+Yc14XQZhBQFgl+tpviSnE+E22lLC+tHGp2fGHfTjag5PFOoM+7DXn
XiWb/tQdJWCXfO2EfQfGtsN/GJ3jEcKPxYqd0DKcgP/ERCLoSOtREaS0ePusb1GOrcp9/cOBFzYo
cz2QEEIjnikOXQ3mJJzQqG8CvVHf5zhWME5y+RHTGUtERJE1nQdc50zQJd5KDuij5oRgKMnPYBnd
mfFN3EM7qzjakjNFl7F4hBqM1FYs1TTYXMDWEcl/N7xDD0odXQq1kkA+RzKnUhQik9+c4XA+hdiM
CcdxNwQD/5vIWiyZnmMePuXAmvMXPu+UZPGEWKbrirlWYDZKKQs3tEgl2cxLtzkSYaPyVT83a5w5
UCJx2uiLc17F7p2vKnJ4kcMP9elopA8iqNfsIYDFIr0xMK88Xibx3BbyLi4q/z68bHYyKTP7jKkL
dTpBAdA7KwQCmzMwYXsNHm21CXQeFtpkn4f8li77Cea0X7eZmg++HxI1WnmYOwkSWIiTUM9c8GmV
0y7VaRbGGAgx152bb9iufm5z+GZ2UxJVPexQlAVg6glTXQ+wjT/VCyl4j8+7znz3XiBiLBT6eH00
rXcln56szXl1hK41CRXXxNzjAjsgng9ZUojUyFWAaEQbBVrU+fyf4YQH53515c3Lkt4axcL7CZAd
GjV3ivMSDo8zEGG4nEArQ22iwLUyprIsWYRnfHJVZyaZ4lBDRbp9NJX57qRcKyGd90DLmhj6X22w
x7jk55kRG0eQ/wtL6+mMrKv1uZtdM0LMn41twJlvfUKhYM57r40CEp/fIHwyF1A6ABJ+tqHd5Wv3
8Vkl9q6fbyRXeHsAuarhkWaAAlhc6Pk4/+EuK9YDBoKT1DwkornGOgxb+BbI+ZcOmSyQSmjd56LK
hM2FKGQSRFgKHEDhCFbyEVHbPNlxbKwFlg3DoeE46Hwv8GOKkTi/XCK1fm8dyXTLgdNHL3smsbDT
hawPCIRkX1fRdzYpNqXBdkI6nFRngK424wOYhil6kFXnzlxIpD4eg2Mq8otjIMG5VAtM/1A2Cqiy
hvfeFfbK8PSWQJ6AesDTt3CEfP808A1Qsps96OvIoCKpF0/IfEB4kQjLRBH39LodYMCpqGSbFK6p
vMJsuwXb+7cz8lgKMzgqQcoGyhr/CAtnwOxt/Gfcu2fG77GoXT/xEge/budyVnScJU3l/iX2/z5D
YukAKaL4M66eqUa77lrtZ0l5HIEATGZTx7yEIZK8oyd7dvMMJRtDX93o1dLyZM7eYAw8uC6yPZEY
P2tTZ6PyCJpi/jJ5CTiw/Svzqrjxbo5BgMpA0NxWQue6uWz3p4exbwc87wliqQ8xBMPEhnR1/8Yx
sYJIO0UD0rlSBQdBqX7qptnECrHWuWb3QWp5oMKMjAYAiFPi9bC5Ixi9A4lwkDQ0WOZ29myKeBii
n4deIC7qqKP34cfB+7xJLGRiUViRzCAx/HATYGN5W738d+SDcBqBqc5yE/UoXME9WXzq/3cc/ctt
01nkMzBf8vuiJeXFHXr4Od/SIxdS4eb8ceD5m4mjRihdohhmUcpag2JLe+2Ium8+y8PO1FcQ8wB0
zQNx46COQbY2/5ZHIk/Wwau/3cA3eOR7rzFZPIiMar2Cyhcza2mNt+vrZgOEaybjS8pVjtTfsXge
yjIOol13+vAokf23Cd73reUQQ/bD5mAp/NP8Jzrpp6uhPF4NPGLlirUh7IVmajQBsAcUs4qaYBBT
6zWBWmrqSeLUEUI1TEau2JqbBdmnjDbIGukB6OfQd33FcV39W/HB3nnbmcKiqbVVmt9bIS7yFnl8
7EjA/NblCzj0LUAaTqrDV5NWGxoYKNWA14Gu3kmY3axOU+kh6oCqlNjYxJZf+HWiGq2yU71E5xXH
KYGZACJdUv2RlcvS9X7O+aO8W+Nh1lSRq8PUMlfLpB6datp4aKHtmHoSn99eBI4q4+jAHIelvpSf
wBxYOoIu97cT5NEbya/OO7nYSQaC/RcrC+r5YN52CYxUUcahSFvVSjzpqblMrA8B0n1znQFzl79o
OLP+0CMz+TO9MU8/gtcwb6h17Qt1f0wnB0tkUCs6NiMkSbTlvFnLjHJKabh2/5bBdA/pCp67fpNz
UTOVk/81+K1Ulep2NYXU249ihN1XJmh2S4weuA+DPbPvsOcx9dmwJo3XQkOv+vOXqt8/Kw6eUlsR
fyd19tDmqNQ56Pe+/eAiGGCdkqhwRLGYtya8hDsSYnabsdI8Ni4P6QR1MrKP0wfjjkYtJMfaokNT
2+ToDOmyaCnm4aWwiiay9gY8R7cXKvhN/RM2xviYttqzgbxEvdxBOZsMQfniPxOLqJzdUlN3V4Wh
BWJfcdUrfNR7jCgYxlz0H37z4IGDGKT717cb8wAoMuyY9Hn8K6OcwG/Wmfx7i/tMsmK8w54dG+ks
p+k4B+gbbnPnUEOvgNuPXGUMOnYV+jUdshu7ORucX5AS0HKS258a8iKJIICET2m8c7kKDio7SbWj
kws4J115e801tbdFdgqngX71z2ZKjZKeDoDSPa0lMpLKYn8YthSshLN8MKLAN9WEKxBjQR1aT8CC
3YHJ7+k3WAO5SqwnsMTmQLlvTN3tmabZSHUY5pohpuS7PJvYw7FfbG792m9xd/VYHgyDFxQ+6/f8
QbQwPA6wfzEYZ/KAkfoJEzk+ohfCi5OQ5Bi8a8e8atQtz9mk7lzuN5SQtDql23aTpJp/SWVEQ731
88yUJHorgEoNQuOBGFbeSRInBx5SxXDzmwVb+OHXPSnZ5kk6pIZw7MI/QZOv3YUKqHdZ2j6dkV0/
4U77CZyFNUKFibavYPcfqkeOkFOg+BQKQB9R3hllU1wa7e314arQzedwxgUKKNSYPy+YEC/GEhSV
uxio4Q6rEcZVelzgVLS5MljGXc0iMcN5+fjzdWffB3oAfE/z8HEL+w/RoQqWgoLYqJ3hD7q0UahP
7BCSQgoEHUVTfqO+hUf6OtAqTw7gBhEaC/tD3P+kf4pfdWtyD+vM9fiTsq5wsVejwo28/VXjRNt7
b/wo3oDdeednw0jR/c0pmSSHt2WczlBfr14XQ2/xo0Yf1+uNmi4t0YcC8/scAM7C5O2NzboP8HOt
vm+jB6tuTly3XFQNwH5v/Os42VGmE1x9EBWM/BjQwXMX0okNaKWpaq/7I1HoQQt6xM6u5THqlThJ
mYJQ8DKDGTo2cEQ4EqRXXpn3tkbRHrl9gdcqOAXTb+hNEnaBoQJpcquFE3/JzFR0lgAAFKBEYt3d
Zv2rKR422bh/HcjqGnGbOXo0HOAd0si1BAjcO5evYv1jO+9Y0dX7CWsi03pfBg9liTPU39BQ/bHk
QidzxmczWhchOH8aTJqCON4+/I2FnxBI9RwQF0TZDGOzcjR5/RtfLeiOlncsKalC3ATDLKAx2yrd
3Ete1cYxQ6upg3sHNy0jANMcHPgtpoRPAWhDPNCx4NJeA9GV5BvOURDJvO/qv1NVGUxqnY5AJCJ2
6NhUK81aZF3TLftHZ0Xip4QtvIgPCrV0tCHmlnHG3BVwMSUF3gfw0w0lcP716O2xyvIwUQQNzIcR
OM8yaWll+JB98pCDMrmizJClGUbYKu1ZOp69ZSU7LPfkely0hdXla7XKpaDX93m1LpovMxV0qlWE
wGLwOlK+UspuIKXCF10ZobNWxzvuu++LHFqK8GY7PNsv8ilOW7z6hexgLpDDN701Ug5S/NnmfhTn
M3VjUPFlXIALIIm44y/QNpYi9rIw0PhWzds9tqcULHxDrL22IBYcrfBhcUR329LcSP0FZkLFmxUQ
KKt4sCb0ntJi5Tze+WKX/NcV9JRux0ZpXB/L2R8zkXZtVxXgRmrbzDCPv7zqiQPilRKIivLUg9hp
hjhbIBdG7pbLfyru5CgTekvQRmRNJ2YOUSccGMdZOIRwX+QMK1E023bZMOi69FNdHkuIFxSgOCah
/kAXBeBmmIqXsV5nbcImuBTE7gUxUR3DzAcYbzS9in1yu97wtp1WuHkIQmvSoQ10AH2OXK/2b4s0
r4fV64BClFPAjK+1Gq7KdAg/kfDBzZ8cw7rVC2Ei8T287QsxzJXueGZ9eqti2pPoD3uQaIfCIrv9
NxKr6IXd1rf8Ayntu717tQE3/Q96jZJCLIcTQHz3F0BV4MophpksJNe35NzDZKlNzRWC4/oo2I4f
lu85YPaRphEIE/W1b1TOMCYigrHB6xjeo599AlvjLl2N58Ax3mHrFB7LgvGfOrVf7IubE+/Pmt3R
vzmf469DTinGtqYwj6w5KOGQv35ADUGKiHOixx4iZPIBQf2567vDQomjQg/y34qQiFPQ/vOCvaCS
Nfj/58ci+Vv9j3BNVvC0KnKrA7ZDveu2ItiUOSSFHAinM1kM0y8xEIgp2j+ruQSn8sfe5wKeF+1m
MZG9/2YZSezQNqJNyY2Jvcdpjt41cbFS9AoSheMVdeinGQ4zeJTZ9OzPYC48zmxohChp5hNV2pAG
yBJvV/t2De3So/7ek7+hph3D+sapU1o9JANo2pAYuDNOFjdqvrBoD1nHJS1r/4nSE9FHSEZSoh5E
zxHXbrwnDJpGsti5ItzcQ0el4p/wOagF3d2tVC7iE3Dyhftm2qKpNAKPxE28FDp17/yjyTP4zgSu
578X/8lGDTYfMlvYf8/F2Xfb3uiCUVNsOJpf1AVw/M5bnftk2ZeNoSxnH+ansC1/BHQLbQrZAd3n
0Fs/RZOv8MSFdBUYnozI38Kuf1QRAzblpI/hhATXliMdOq6s4ecoyS8mIAr5S5j+chfRIkyD20Go
KyHl9CW+/lmviDWPsPGJG6GZawAe/Dhzkvoi9ExFvsOQrpjkPu3oUNZE/lYkgw5T4dai26tqN/IK
Sjeo9rJ3lD7ixkeWJPGp9iFJZH0VRZdxE6TpptsYPWyvmgAxmSuNwadTaYj6aTsEekxi9b4IQ8fN
x90VRH09En8+LZpDrkQmGgf+FC4RAJLTyCH4PD6b+c8zQu6EOXUA+2ibAx3tUoscjcaAcWujaF0c
8oTCh+Yv6QJfJBXlu8LBwk93hh2zLtRz5LUdIEdeel5B2emaT+S5Y4Lea3n7XBXDsdxAbBoL+VRG
5izCeTYqgzN2Rhzj26Nl1+zWjw9GCjTZjphs1dCl2gpBPDyXSvdcklb/vd9EBHc3aByRoYAV4bsu
8dPP40HzQfCBxxElL0dHcxn3fXUv8cJ8uQxl90raaqiYRku1sSjES6F/hRhfYRXt+rJcKcAVRmcr
RF7VycfkEo8lW87cqZTtZSCZXIfyCu7qdd/2S2fzX1L1d1ttymET1BXUsoFqCbQHedY997Y+Ef4R
5HylsVpFWCgJNf59MO0liR1ubgU/FJePdcU1c3YLdVxXYxnb228hmQ8eEtO/4QlxXTOiSvC1flSB
PT6mefmZ4dbwz2A0ZAQ+RweSW8Fe9LFXQwdkoMeNoKXce/Vrv3pkrXVPyffNDKZf21kVeb9Lo3CH
o5MVvOt8TGZGSG6RZgTueTWWlT4nkxPX2b8yDoxclMGNlgaE0vuHjzYkyoGodJlIZduPiv+kG0t1
0b82KijZSrf6J0bSfXnCl8C+PB0Xj4LqrgMG6kJzwGuq8wW4vuv1qM4OsgZYHhXWbmQrwLQeu/py
cvcMWDXupUGSRfD4Eevs8MPTYnHf8q5mkV+xrOeTY70K7cX4g2c4Lht3KTZyFbGn0M4MM9UeHyS8
gPCREMJlVlttXgthrV6ROzvuZ4gNTt5EdR23ND4FlR4kwgQcRW6nQvqfR5iKWh2Wr6cfLN9/icKA
fvMl5PU1PMkJ2lkFJjxBhcoPwstKLfqVE6fmelBtznCrazB4UwQ+8V2r5f/hPi1uLmNoKkbS4r/2
REEGUnI+m4YdsTSsWsuiO/2g05nQOqvd39JHScetnG9e38WfW2RSqBDEM2LIj1/rc101aphFii96
qajgp0Md2N+GILmx8CyhYKOYuNBxINthHjcLJJ7dNjuid6TiL7lH7XPt4P0vIHoHshweKZdmgjtX
o5ZQONuiPKUfpqFUvmk5WOh7LXYlEXux0yif/cDbRY6B/HuHMa2mZKlaRxA5uGwEdnAqjephK4Qu
NEVZB47qyDX4MU+PcbcSC2dA+x2zldXqeGjpRtHQfSFhdj5dlOf0LcPrxVhzmS8ymnvJbrXI+ys4
io4+06yyvghx+0zY+h50Lrilp20YSuty1kX1NqrAB/J7ejmwLwjVzek2zoTbnpLu5LBt/9XODydd
H4oTy/AXYVpyC6CdJBWe8/qwMWhXetcu5Es+kyID8zvfL4+V/GxF6FkBZOYNwNoGXEZcML52sR+/
WEtDZ+g4AoesFzBJ6Bd3UYZLt0ZYqH62FtLx4sPjDPToPL+m6BLwexou12Kg+oTP3YKfd/evZ1DU
uMpK4r+64mhirX9hK2wWW4NR2IhlTJpTmcwH0Dm880MRj6ZMR5KKHFrwqNgN5FuPrBSTN7QxcXpK
fnqCAeNmy7XKVGvdbCNyorp+h52TsdZxqN5pCtEsOnGohcOFQ26dIYqYjDJoVq77k1ZiGbRjW1OT
9+QXBVCYeTFYr3GLVKE58gKtycLgWqbU08sIxmxv5Uc8flwHQWxU143Wxh6M0LuYTcvMijJ+4s09
MORh8/iS83BttUt8ot1pwLvRZ8m4IWR6FECTkkFAwjyFyboW0gt07XHkE1bDMHorHObASq/lFIaE
esWvm5mGENm464RE+kWoJ9YHGfsWttgUr9XnV9VKjwv0vwyXbMC7UrQD02yZSSD9S+f3C42xp14i
ibN9Iz09srDi6Savq2nDjgYBGxX6s2XFGQxLDNWH700ZQcVYxpKsosFE3ekkhrVD1jTuYSxkdsNv
S7/K0HyUkqmFs7Rt+Ygq02ctFVS/T0DUE3ZIUQx9hwrXkpW377ILO0ohVqLOZCniT3hvS1KZQ99d
ht1rIEQ6UWL1SEn63Wmlne/wQYlIgbHRsYX73JckbdMpm92E2xr4PpoqhuMNw3mztUJ/43tam0yD
1T1PnBHm5+7kJWnKgyCuQrY2hs+UvLYUcWtEZBZtw5uXnoFEEQmKuB7KZlsB2q2655rMMVCqVaTC
IzkSEOn7B83RJYAbQKV260J7EDBD799s40MzhmPav/+R9w8HDkFij+Hdz6/qlmW0P8uI/Sn2AqCS
f77E8AsW+sTrWnxJhPu+C6GmeOyeFq+BarbP9Ka4OFREkIUwyXtJCV72BMwyqEon4/myilCvCudA
dqVRWKephAncTQD0Mdt0gLasZPmcfVQ5Eo4Q4dQlU++6OarGv2ilcNcNxLzd/vcD8JZB7XMl76Aa
ybEDZ2AWkmVUMK7SLYdd9mR3z92RZtwovbVDhiDqGPtAkRJlkYzXjzkDNnEPQIHyryiLnA2EPwx1
y0A73V7mR4p1RQxcgbEwOSajHogPEFugPWZvfJAKCkxlQEmZtY3idjKW2NzgPaBE7Wmih73pRNxN
1LxNgI3l3hoq8TWlu4W49MRfjMs7GXNqI1lNwlGUdGXKHgL42qzMk7zGdi3VUxgbfwSq7MNnfElU
+R//SMugMDnMDamXgIqL7sf+uscFZwXgcyxGGVtRTFNR3xRnXSsSMSKSOZ7W68PLpcia0NJiuqj+
Ee5gkW+rW7Ge/HLm/WFNxb4mr/rTA8ZfIuxHI4szcz/0Yx4xhkM27rErzkFKXEsLDRhIAsylrqvn
lLlwIZ+hIbMGv578DmGyalbEHGAalJREiGGXFeknwN9yZTAhfBEYD1L2wlifz4R28rIICxKkDuop
YM9yNhEClX8/yF30E7Mp7mFWYb8wDLUcUHvAYQxBTycANKON7jZ8fXbNvmL7L93DbZpNaOGrDv9J
TrH3Ds1KczI6Ul99q+UPcnsZfZ5jfVbrp9nfmkJsQ16IrMMx3ojt2l53djFis1fSBbSMBpNL16hG
9oYqTHeHeB/ZsacjJyD7+9fQfqeYeOnJtbyWcxq7ElA5PNraqeSXk3IN5wmuPyzqdUxngnplt46T
cAhMbAar4lEgB8gCthQ0iUEDx5xPgQBQTJ0zaXnnKNcerpDz8vmDfhVfUPR2+x7IbOSeXKUCRGwU
aN2tUlWq3ds6cZljaAvryHbVWANz2QcX6q0WyQDVDkURvpokkRXAL+GjRXV9tVbk9+lQdqbylMPs
HXgUU0rsITHCMitAj0VqCaznyOBut8bZIpZ0mZrwqvWLzmeE717gxk3tw+u3EeJCljjNlx2HHKS3
orYMyeDYjJWOetWJu0riRlJ/w4MYa8JXK6m69ZvebiQu1x5tXE2iXAuCpjz+o+g94i44cLo9uz7Z
3kmzVZiMDiTvxdoSBBegu5AiHdvzx1TURYfSXmS9th00cZ3NFRqwRjkW2h+T6Z8mtw4/RlkftlGx
cqWqGOW8NfLqC7TarSWd+obfV8CgKM/m+fxBAD1uVTJ+/vvoQaz+qW7SzRM2qR5Kj0aRLMfUaJY4
uRm6JsJe1bX9lrx0s+o53lYGtpoCL46B1k5gwv0hPt09cpQUIfxu1nEppdukcf8w1zlgEEMdCcPe
06L8WEdIBC0gXBdXlth9dd6aJLZb2DfvP66MNjsNSaj2Cgo9m+0YoCpM94XeTq63mf7EFPnVkYUM
UmA7hNIDUXbSoY8GQUDjg475K/hmClLFXMyLCBY0Ha3d5zzymnXiDwlsWxYIafpuRPa95e8EJY4a
cd1jHgbjOlnkXkg9hzI/YE7kOoyh6KPuytG084kY7iFvXFUGEBjPvcXpDy9IYDHugRgUAvokDkkI
qTcOugPrqdN2oI45O4mobbN9k5XuW6JFlS1CiuQySv0PeIvxoR0vNuQJ3NbmuSHrKGw7szF4Okas
botSEdXjzgO6GP3QBXsBFpOI7oNFWNRpwu9lO/F8XKDrm1NQ1rJFwEhehrHUfcW7lpJUTJqb0DmR
PKD659D3jVPVaP/CId5n9R4rwEXxWqiP9lkl5UPqf+rvYvGiDtZWqkHwfVJoRKownITmU0Tgy63F
PGE6D+ajKkIV7LDHtfu1YHmpWNg92B9BGqpnS6dWXSaZqClSI8NkSPXw4rHgqroJDq99dX27qfEI
OTTnNEHE7br3YLeHAaKLmz4Z3AkEMaBD0iUXubcmZQkTJYKlSMTxV+KO23SrHvGtIVgwRgSyVCfS
9tklJyI2snMiIW/la5LILqq2C3J29pk0FT8S5bOYQUgTg4Q3Q5+7pnQKdmOb4E5Oh8VTXeKnERR2
NbGjEr5tBokqL/dFlcmItIB7Ee6x8WCqbmiNBvBIMboHkcnqo3oRY5+6ISqftNrvcY7loh5paKZa
3kcJenyt79SohqjXeXX0uVU7OoB1vd8IjtNIAF6q4hnxFKTUPlGpzuJGakoafgyHTLPWIYeBL+oR
cMitDrSdVo1LUSPA/1oFmRg9eiZGnycvauCYkevJyg/j/okoNCJLVHCqBkYAa085Y3qroUfeSLYe
dtDWkMO/g9NztmeFUSdUZiDqXQPMJqzad1ltrktrlKbEDp/eG/EnxBbwP2AUpiRSbikn70qxiEU4
TgFatkO/Fa2LRQeQ0m+QX7neSTyLn98DXP/ercSsdmD2G19lrhBVQl9n6NA6nyM6zmJAm6BIrvWv
24gJFPxDztVi6IUhODgh0InBQoFsPMWuUtPSjRorSaepJmcyODG3M2fBJE6Nk1qi1dsCZvCbQI3h
i2RCuWZeKyaNGnq2SX0XhLbaLK1Vkg60pF/yo+NSxTVymVfXV+CnD8zPfkAr3ZyysmTg66aGnpKr
+R6GsU3gNtm8TTjUqZZ+9ToI8tNaQya0T82KR9TONXYVhvDhaT00jXNf9ikXC48BYpc5o0OxsVHJ
YF+PEb4G35COAutMHtbJqUHFTgtfRg4+BPHK4wQN7n7Owc8cA3fcnX8G17S4F4niQLiuHPL9je4I
0tvC8TLinb0J4Y9W7hJSqkZLOr8RZ924YTF6vqi49DXVlO3D4KhnKOAh7atPtZ5RItDLYFFRPLBu
mSEvFvWiQxyxor3nIDMKQHSNv1OLDZER/ww96OSnh19DcHXAW87supwpp0Lef5zGVUzesT/7OAbV
BEKwpuSwnPEG9Y7BXbY2UK8YIoZmnPpi1ax2EnSO5KeX81em2jvFuu7FtxJOzHLedIaLjaf9k9xW
kKp4Fv+ptjb6Q0hfOgKOemdnYoJ0ZJulp/xhb2HrbOJmMjDzhVIy+SbdE3NrGHFbj5UomDT+SCuN
AkERZ5UtYiNGUambydpsjFJi9a20WTw9a2YF8/GlrIotTPzAAjB+TwSi6CGTkd90gdnljubr3jye
jDLOc1oR8mM3ErReWolTUqXQW0/n8nvPzt0O77+ynQSU49iXAYBOMRewZLQwC9opQOj/S8IBtlGX
tHBMfkYDZ4j5Pp6ppH3BQZqVFhspITtWPAlLVuMIwcez9lbltY96vhUprW55y6v86HJEO8lwGT8O
hR433TO082S9/BtGblbm3hcYqnB6qyVWj+cGGvGapR4LcOovobkqwrjQ8Ex4ivhs7XAxHGBIWbxZ
acgZgr3Llzd2n5gFX+LxEn5C6UmOgl/DRTMbd1011SCo6O0HJcpbkml/td/YvwP42Y+x6VPIMXm2
tVVfqY/+or2beWCx7DRhjuQvIgLepEYnn4AxX7qE6rZU3xFCJ/ZKrG/0R4ZdqXjPnUp3V/rWI87w
AD9djmTn/4zdKqexu/VtlbfVKMs9OZJteRK++wX1lF6qeq3GRM1AOe911shZ6DiVEcEvO/fmVlko
jQ07+4o6dk/0+aHSWaK23Gp0JD7XUn5xYQEJa+Aa0XKHSI7v7Cey0F0+XP92i2kp70DM5Gqs0ilj
n/pgYJ442tlXlQbguLqnRupAwTpy2mXIqnXMiAgrXujJ+TzDgn89aBVVylSpxEzdWpZGxNoAExlL
dQYhWB2vMIVEhiRHp/+3np3RAEY63Th8rP38zJpFNJ6wPHlkOTfkEUuprIpKg8vSjmw3hfTBSPja
rTR+CppeJoZkErb7T0WCbEjWfcBoOb427+pDxVdS6dMVTrv7ONMzPcwyWRDYOXHiE7wm05I+nOJQ
Hy08VL8dfaOhx3jf/tB6HVaLjm49/Qll5+he+L8GMqGz66MnlhsFFssMjgTFoOkR05xZwcJnSVCW
+ZPhpmU2fqxL04Jll6Cr8gQF1JJ+JaOlsgq2hrJzjFX4yQ793Ye7KU87qtD/G0tMh+o+CjPnvA6l
WtClJBhbEVM3zSm3YzIOjv8gxRFbVybOVx4CuH8A+DCQTEJFdf7VB4eY0X71+w8k7uUH2CnLmZlV
pE5oEFAnOgHxi+hqe/9clkWqQ/w1sgWmg1KhwI9fYnyxlgb4HUlvMkhonH+S59vUbVoVkVDbwyyy
mxGY9CRLUB4Bef5RPnVE6enRQKSsGAmMrXGTU7dEkfH5EgaR91DlEOqvfBsTmk7H9ea8cngyxWq6
wSfLkZv+0iq4PznvGkCs6jG0XZlds9I7+6LusJNLtk9hn1q29pfGscnSRg7nwAZipQ0DXEQXboCR
c/8ajFJTcHo2hQ2pIxsSCS46yH0gPKPaU9TQA7I2wXbW59b1LZPtHxLLw3yKK4QIpitZKIr7fn7e
y4PSIrA+7cu8oI0/9ZYWgZkTcsqqya9ggqewmhmBeiEk4JVuTi5O237eHaYAGh3u+9wi5pt26l8D
2t5GhlCvqvQlh8x0PeygAt5ZzB7chcIOUBie/yJ6z/xHEYZCaZNjNdFtac7JuG+qxAPgtQggGZII
zZW24rZXG5L2B9tf4eUgQqx29dhzHdMrSfSCJiJS6kB5MjVtIvWtm/CvZwsNp29PLbCgzHx9Z80p
hH2T4AvDx6zZV2Kz9P64dqm3yoMEEZlRnAoxYSwI5DgbyFtrfMsWTjZOGMxBcjLkiwsZTt0Pwjxr
rLHEK3YqiqGXbfXlW1119h4PIA3Yipb59ah08dFYODCvE4+ILm+6bknUPDe6drafPzFrh8w0YLsa
UNpZ5/jQUqgmOS1/C5pffqIDuWPD/ETH+Ybt/rDlojQxHlSEXv06UxISQnVngNZxD7tj78cKOrrV
unOdQs0P7QIpAOSKTXefVRoPJGu6GT/TXrpRJNY6fAFPpZGsJE4MCk8NvJ2onLG7JiPy1GfnXOIS
mR8FbrvLkTRIqJd7Md1pOvxOtK8cqhAtHGBozGxy3kTkt5BI76CgiIFRNXHPZgFkrvDQ/9YV43t/
ZvcHwM6mSCS5nNDxXL2+M10V8dKz80Oevc46ynWjfzgbZqpvB054ikO28CREL+qaltDdrvm0XMSZ
N7+7IdgWnH5eoatVMWm0kUbksQgyMRjOntq8twgFiiZgtz0w0jWh29XOxnsZmn9hiwRA9S/ll6wm
TiMmrGkG/EmOp6LgptcmtaPnnlhANVQqqi7u2jdJXeGE7G5n2KiXQ/AuYyWWYPyuVhNbUE4IkXiq
7y9C/SpmOAXjz985b7/gT//WoVynYf6fDuCvz0MavNRkFNxWRnP7u/JICBxG28WMsDj3ULzrKrdl
CbDy9EZoik+S7paxJA/xw26nZ1Mp7u6CRn7CGx1gjbU9YlIW9KyMCiojdb1PljJLK1PmuOlBYxuV
mx1jD/WYt++YY2YzBnmyuQ0G8/oBdz/0yeatub1Ayx3wrXWTBrMMaPwxaX2f1hdLRu/SX6Ndkxv1
13F1F25LzOrRZ8SchfFhSv18V2yjFg37Z1QA8LrMKBZf/LpqGua0ndmM0ticZzkpUcd/ABs8EZeJ
3MtvSX9QIGZRdHomhX/5XO1qYeZMFadTkTG8vxeh4XBGUDakWh2SEtGcIP3GYDvRpMom0/++hl4j
AoIGfmJg/X4XKZoV+si/epx8ls16H4iIwecR3SAYncHp5VRAKL6b35a/o2LLj/Eh8LPiVvMoH/jz
Suo/J5Rek59RNU6MOHcukrVTwUwoIzUXJlCUxsOMaOaR69NxP2W+RBNkRjABTHsZkffCTsc7N7ui
TtdUhj1z7s9HyRsfCbQKcbx3PXkVAmDxwOb5OzqXsQdm8LwTAmI/mFEwsSTsKFTK5BOzbIFP3b6I
2pTpjX7rGSE7KNq7HAzSE83D7SNzN3JOh9jLbMNBdj2NCeE6bsFwO1IU/GgD1jsX+mPhHR2/QHFA
ja8JBOkCeb8KDGgT+wzbmFbH9LMQnE5BLrH/rRFDt2suaHfB8OmErlFdYj5Kx6skL3TGiL9D4E7F
nOMjcNHvGsHU1jfasISrZN6vzf3U+tC9vljnHhwPhfF6H7ax6nhaLm+lTvUtC5Tfgcu4mgxs1AM8
4BSHOBs4il7+S7lm3cQ7fs24612J5iju0TCHCZ5LQO6yd/O8BCGSLJRLql59AkK3bpSIvcZxDFMq
z7yvNQULpIiVpeLOejJNHXiBUkrO6vcrlMOMQ8XjYLTrGnRZeBUckIjTe01S/+7Tbj9QCniYf9P7
VlomvzxRTxRjOABpR/l20ARstuRIJYJlLAXBDjtUtvrFacGK7Yn/Hf03kT2yqmbLtIAFvuLNkwkp
cNcA4J23mjb1J0lFCm0bpVeE8Su4xE3ExEfNcBuk/T8O5uxNGJLgiSeiC5Y5f62hS7RhTWzuhycg
jkU1qG4jgzCvwdhdAVewXyfbdEMEM9pzBX7Lnyixw842MEIySj2J5NKW3WNwDZAI9zhJVb5hwByx
iA1c3d9g8tl829h5QkKwUFmAldWBwUJBiUeVecRt4iwHtgkptfplQLb065A+pj8C86+hwx5Fw2Bw
pf2hCB/VyBopju1wMlN1Irm4e5LzOXvTvUE2roE1x6TQgQqD683Swjk4maxSgqzsehB0ZHHfwBJL
TIAHMlwGUS1eIS8VUAlJ49en1OnKbrJTRZCsdrve9EvzQPCMmzKyYIQKDuRy7yWLy43TbpCQ3iEY
HvUc4BiskoyxlTm8Tcwf4l2lLWA8LH9Ee2k4tOL0Hgaz4E/Sqls3psHgMb0FYu0MqNAqZWaf0cGW
VQP9QRXX1f25zp3AX4ixpZrdnyFQzC83HCceKcIaEHdclWrXGDR4zo+f7FTGv6dDTT0EOuZZtCE0
9FxXDD07WrzmSt5VawZ3fwTYPwziar4y7kiG4e4U2+Fvc9cFd8krcy92LT3iDBNXGPTV5fCNKjTx
HJBwSW32uh9dFz16DkCTTnnvtkRgE6e3ch77kjFE7nE1xn2dJrPDHPWIkGmqRtbM++BIz6tsBEt7
HhJPEbqUr6einiSC4S9O5jHS9BhU2hS5iYBxKvGXxVYXUWhFn8XIh28L7dp/zDZPvlFkisXBgQb0
vZfG+SybEotQ4tEUgG76a+uetQosqsRa/reFhCuy0/rlvtbwBwrWwB17B8NdgUkus6gEmzjt9UeO
UUXzDe/et+w0+XT5sKL6976CiKXyjX0PvONOHDdgi5gYcafaVox0qzWkZOJy5n8FH8Ck+xrG8dpI
upl7cZ4S7Fggw7M5q4fEAD+sU357/abo7XgpfXY4qIW0VAxYGnoJuh+4GThDgQktYRPJyPC/4gzX
jfZHJDIxN7zGZmDEHZYB2NBRIUNJdLQqSUgKrIqjyJIvKbHi9fD28KbrsmDvIVzrcEieFDeuxz0q
5Oj4j7nVF/rAcgAeEbRBh5QBLbJqo5wWrwL++f6I0H4yYiZ8mqQ3LPjLIxfrnzBvhBmCYFHVnxXz
7aHBkmo3zMSxnqvvAfT234QCIHiZhTsv/CtsL44zQY2C6g2UPaOjirx8CBLFMNerfx3Aqu5uMIrR
DIZ3qPm9QITjK9PddZm8m7xwe5ViKme5NbqPdAMnMYsEdxxgdsupJfEAM+m3StJfAzfArbHJ8azJ
puX/7s0jwt2d7P+oCV0AR3Eeoqpv0IjLn4yzMCT4NV9L8fjuEqJ10Fo+PUFWj4J6ftSgr2KYBnu5
/E7oJPkmbSDco3d8Hq1m6wlZEoWWKKZOh3l2JHcvE7Fib/BuqVr2kXit+Y1vu2h57H+jCW6qMAyT
1BqGQVnzT+HNV4VIvoHhAMK+Fcezd33ovsZiXCJdQWtN5TRqokevT7ES74lcfd9Ri1T2/KOahx72
mp+eBNvigI0qv+HK3rPmbjpDZsy/XowiWXjkhVMgZ8bT/maoiQuBpFs+ABTtkrjk68gAyk5NOCm2
xd2K8t6hr8ZNgcGKXaQ0qYJEV3Gk0v9PtCKl7e7E8qUzX+bp3WfhwpT8Qy0u/TM4/WKdfuqWZkds
jki+W8MzKd6cs9t9RVlK3l3OWV+mZizYYlkcM97Omuw+mI70/2cj+HjY5gYpuhwV4hP5vHaLQtVS
hXe/UkjaaGtQVx2J9TZ4i2RWff3fqGm6lGaCKAIw6ESb9czLceptyNra+OOq9Y9oJVxzq2xe9PoQ
vYDeclENCrG4eXmZBIbARM4VVEfefYrQy+EHAhdW4sdQnUNaK/nemvA6gWqgczXNLwD5AEmz9Wuw
g9+lPbb2ptPhRWFEYfFRS4N06JO7+MYmUUdoHJiUQoZMidOElKEPQS+DBv6rFYX0362SiY5KjCnr
PrUifvksL6Vxy+UYjfIf5+Lyk4a4K5SAzDE6ij9TtB1Hdc1KJCV9WHe/76U2fxXMyXPEp0Qj5Zu6
iHr75RrMmaPXxiLI0AuWp8EoXuUjdJIlhN1HShK2WJXu7d8aVgpvH5fdN3Y2Ylx0Fm05Zcbss1oS
3zkH4O1Bwg07Aum0tHXn0scSYWieZ0N9vRoPr4Bn18p2oLMviYE4gDkOjY4TPBje58kiSLHI/R8v
FkbwcLU698PYWdcXrIQJKk1i9AEY8L96+ULbem+7cjP15q2Hc+FiH5ECb5KUVgo5TPGmoC8ygCol
RIJ8MwqjDXMXlOMQ/jNhHgnosFn131JKXGRUQ7I1z/7SrBll6BW4FWaGHkGwv+0vn9uydtZeJ0OZ
oQQH+I9vqGXq7sUWFUzSQSyea6HORLsELK4kPKAn/AWqhB3yjjDtGRF6nh20N1wN5BtQLh5ND5CT
REhaM1scRiTB5yKXdsAu47b0OHE0KtZBc9im3mO6cqypOGJUB8+ALm118dECoOfUVMsNsWVyWVs8
EPxCmyjzjGJ0INZAH7yhOi++/nqqwEFKmB8zmLPgIvAnEii2SexHRgeWhl/ko6bUW52CvM8BFmQj
l+HKPsaNSar3O7+6SirxUl2kPqwbi/OZi3whrHqIRh+kRc4rtPfIWRiFc+RefkllFLVAiHtdEBYL
fCCyH7JkIl1SJMhApEJoAWuwhv2+WHV6QTHfP/xOf4Ixb2ZTPg7zIDY7NhTlOo2JOWm4171tHhuE
vXjl52hVG9pMY3+yUTPKIT0Zmw/IMsy0LerrzfDggKuU0q8mcQiI1niB4diIXkux/tpKeVx/oFe6
X6q86O0hHBhcnyT1ylAXaycFsjBmHhOdJSdhxTx5a/j7I3otok/UN8HOyyYoXwnRcH1SgfQQdSkR
Oop/lgLGUQcyXK94Lv3Vg0ryO+T+6rZL1TI+GELMKy8/JRdouugfSlJ0nQx7J+9JtCeBQRBzJfbp
lstL4c5vfIhky72LD/Aqd+uVB14DN/XZEKt60au8AMxOHTpP6LPtCH6eldJjbdSM80I/D+FDiEqR
dT0mDRQfWze8ZGDgQ+ewpcqUBhFhpT0N+UHjSMBQaXKiS9QGDAeVC/ypHVELS2imicAZx4JHciso
GgYtGAesfbxrfgi8xq2XqtfXkvnZFKWnR+Ct+vLNDKgzfghXU4sOr/b7LSP3BS65xskkx96iqYiO
z802ejoGtCko5yzLeV25x+F/w1elpna9zwG4VMPdU5HbXwTuGmVKSlhhRRI4zU9Lju5iJATym/Cy
/tF+TN47p14Amauvqq5UJu1ndlLgnvCu1tnUBrfmo86hGzV86JMXwhQE7DQI3NCaMEFo35x5kcW5
xcsfOjBaM91vN4Y4AQnkVUuW7ht/wdbMhzduFNSJ/08zCz1FGq6/GWwwYHS75Wn8Fkqj/mA5LtIh
Nrv3gtpbvP2hjm9anm4GCBiCLtwYjQHgbPJwewA2lFCwoSEQA2q3uoTOXnnrXD3Oa7cq0BCdeW7F
FjTxmLYsdXNVKVpWguBWXqz6pdZWu2Quy6sWwBkCzjyrx6IHumpJ10+zd4gEUeQyuH/6tKI8kCVz
W23k20j7MvCEDGoEcIrHGVd9a7uoRQTMV91KGeR43jxLpomRADZoddw3/f9umJ3OnLsBK3yvj0tf
jPjGm5gCFnv4J7YRFblXwnvpgNvJWnf2WJnlkwN1tucxQ30st5XRHdZJziKyhhp0WtomEhWZTY7p
EnYGkrGXI1bGOlobSCXCObeM2zV+V1rLBHS3phJOfZlYVHf4r72IFxIDp9VffQKxNrefSZ1qqrlQ
Y6mpF08uZNVhkoBSSdgjwUEjdgnE17DlKVDOtw+eRXjLnf/a4CLZrX7vJ02iRkN3Y6O+/kA2MX31
Msovr6HvxTnL73Lr59ULF9UiPyL2XWsDuIixoRCDgc+9f3plWe47WdQz4dXOxIVg7gvEWGOlufX6
aDRoxZU6y96H0Kk+vHwq7TSOm74e/PlO4vVZsXUMIyNN+LI9GDEORdD3yE8dpB6DMxOWQwDSoSEo
8huXUhlvLWS+OgnHfnGUw4l66Gpgz47pAQsWAfiBWHqU+Xxu+0ZQFDFUttDHzhfyDrItMHRmBWHx
a+GLhQhOGnu9+BTxvkexEP/P8p+GM1oBwOyaMhT0wukf8tNRKC/LZbxsJHpQTyg7H4QOJft/TmNo
dmOEAHWncQ2ZT15J02lbaFASGWlonzLQGVgp04dZ5QfwkaFPIfoPsA7C8Ug01abHUFFDqv1WkiNh
G1WS0MledsyaQFlKX6LVbZm5dpA4VRtP06s3DP2cyWNv2J1L+2vo+gYUy68+TivztMS3BOOXh+uJ
RHL3Xz2pGvcqE4xYiGS0s67UAbOQTE3LeywaVjG2inhxDldkuHoM5/DeubLeboeSp/ULJnmzV2Ww
Ie7Ow/BOhNtOPJ+XM4EjJRsL35kHpG2ELY/nsS9Xjzwj1v4RnFzKpwle6uy7DYiOq01DuP3FCUCD
ghu2d7MKIdm19teaPcs/wHTSb6aUwAk3pIiS5JNV5799DO1CIxbsbDeDJVe4wT2NZWwc7JMJPXB6
OcRLSIpqX3Rd9Wtbfg3lGnF/jaXM+0hnkK//7C3Frq1IWwOu4MH2ZBnHm1PHZiJkEvORunCwm2Vt
dyaSofpkM2tNUfwExY/JTCi7HmNvHBIMpT2wZGMfpO0KS73xqu0H7huKBENHuNKFwuuKNbIIbcTl
iviuBJakRZhDdpIUD54vYxshD3bAyp5lr6Wp1TxyebREbMiPQjHcKL43tJIPJ+OymLv7C2RJBJOT
ZuxhmlZQpjMqcuMHJ6SibpdThx02Po2nsvvudtXkoQHstYj80PmXa1zIzWIKfXEUukinsmPOk+z1
hq7RgR4mt6DuJUmZOOeWFGX3/dO5yO+jWSCDDq8qoD9mgzPwP6OvXO4Lz2sdURZQJW5ewy9ScT59
Uno9/7NBLEoAwKGjZTyrD/PpLykzzM+1YrhHkXhlH1zbpNjhJpGp0UzbiNpKc3TJ6ewMhigcQ3BK
QTZ12jDOWBLFiv0CYQaOfAuTHOO+gDLzN4H+tlKd31eU98UAX1zsmjLBX9XGTisYDNAyGQ0QE1RR
7eBcV8BHOQE3VjsD/lZntkHVRfJSh7TKyCvGZdRNTe9GQNGql7NVCExrW50ZL48HhTjNxGhkrl7W
oWhoaMmos0koqQG6JU0UFHi52zqrd/AXr8uQT3uxA82RkGcEh+KNa85VbAlLkUTi+9zlnlWTuVjD
m9QCdbvTO5mt4JkRKcUgjS3OpB82CBD0YxZrVk42YnN2GVDWQrqgFq8RG4Pua3Yb4rjvnt2JUx6i
ZXeMaqG+mm7mkPpLL18CaWQEkFz0TJLAnhh6tpydplXfBysAq9wVe4sJ/xOxQVS6BrQI/Q9a6S4R
DcxfwICP0wyqdPI8MqHQgMGBDeV6kyMSkrAOl80R+2uFpCfE+duAqXqEDwwyuUO0Rl45KBwUyteX
YS89SGXN8EendWk6XrBX3mSc+R1Safmg8ut7b8rcLwTSussta7pAOgaAEeAT7VIn3AH7b4E+i3oa
ttjvDLDsWn1RNtQyBHaw5QJMzngwbKu4RSKDpZYg3IPQybvvm/SBewM6xwlb5e06HPV43/76w+pq
v5DxQjmoKkY0qpgdGgrvfudu7Bfu6imRXLqB7SYzyOh0YrMtZ5HhZ0Y5K7oW7MjwqKtc86gxnLuF
7deHlbZgo/7KO77KDld58Izw6VCkS14WFN0ucM46/YDV9d4/G8kQcpYu+X/h1gNIoPrrOygHx9yE
8q7k9a6UVmTy+a7RqB2oZ1cI/wsL+n7ACDGBHXE+R5gRoE9J/lNLqm4IJmga6SSa9aBpDECQHDTf
tHq/Z9aY/DT98wOxe73hpbpXgh5pmzVYxz32wU2ZKewtQSbQG8QD5htDukpaoTteJMrrOa3RaZX+
Aigq3+VIhdzlrgTZfc1VUf01Du5/Yc6/VsBV7Mh9iAqIAZ2D8nyhe2+09An5WgVjqVkw+gge0ByC
nhCKrstPqUTGvPdCu0Pc6VGxOjlUjwOBpueB5jS6x4OXoIohhAcI2298S2McCIr7FvS0dId6g/Yr
0EM92YbiUQO4+2IleYJaguyEGmlNkboyJHrksUuKKmSXmZOxM1dlCHx1+/xMqlfHdUU5aN1suK6S
/E9RgRMEjnXtwd3BBeLjIx2WVAPnuTpRXqqTcfTm82hZz9ooL3vANhCxOvUAmokaYtjrNnEoL+Dz
De1BqgLQ8GJWHJ23aGvFZzkieZi7kSMZ0snxxZ/vmzCuBOnmTDi9oR9EMrJOkRWFTYwzK5gUXRdC
5/9AkPauTFcAN8n4MfmzgcrULO2xsgqiNbQ9FoR8n5/I+TITwTspMZ8DSZLCNiKZm8rz/lyPxIlp
ZbY8hY0waMloKespb5/s9GJyPV+gffPpKB2jVxGuLjfGSxgVxDkaHwibTO/3GiXvxGhQjCtWFgHt
QmZLfyyFmP2+hzGFHFUZO23FI8yvJCXbZPjKDA9Urgho9m3aSkp0XEygKjkhs6fvZVhTyGPomWG2
fRk10WJw153E3H8YTk5vghH26J1YVFEReNzuzXytVT/ubeYiUIp40KC41GfTzJGLywRemfWlP9Nv
U4zvbCMVHfVC44T/oR5DkV6oqYJQToOwUVajNylQv4/1faaVS3iLa0IkXth8ZmXOJr3tHuE6G7yD
wl6gAbHrT0sF45MfI84CyCyh98cpB/NA/5ZfSqVCXjfcl8a+oe1L4LWU7oFR+d7+sUCb8rYsRkXu
81aVpt5Mmkxbbd3+wmo2nKa9BHP85o3YTYfUlk4XCpNfltYYbtPStoyE4wJlr67WZ8JOdRrKHbO1
5ljy/6dgATRkrDYFR96nZFpdnztGBBVNqNRZ2ey7aiq/Jc8cbrKDSZvO1nIRiPMnpaA8nMgYc2XI
TFdR+ZWjBiXpS/PPfPCBLL2B708Pwn2Mq+uhb3Mi4OngcUDw8urZXKZ1IoUZuIxAdU5cP7MERRsH
RtT5Xp9yibPHMMpYkbo6iyYcPdHZRPw7RjfAFTV9RMA+2Pk8stsPXKuOXxJlQy34I/eJ7nlYF/nv
oxhJ3wgXVhsUqxK/BVbr3zC6jE2siuLsHcimgG0mNy4HtD0TYswMaN/64WzyFWWcxUIYipF19SsE
Cf2mPhQjdBl/QVVXCSunpDYfGq1HaA8j4asBm3mkPh1Ht08CBdKjh0ktmvX/BeuJyS89FS2QGBDH
DCMiw9AJcXynikQun5C7SnbKZz2FEt60laWUbYJZ+R6lvt9yj7/VC0AytU+GYxANPE+90ayJozPh
yLKMv5knUASbDIM2a5BORsq7/kRjzIZwRxq0Pn31HDTR69KVyO52Q6ayE4kbOKoClJp4I6lBKMhK
bYiV5avtcDBM7hJxjAF9HYTEcK7Y8aQMZYMpce4JQfIAp4/8y3w93EKyUTfLfpRU/+ifvXQTpyup
Hfh7aQLKeaeOVXhYy3gcFOAiZ7TfpnFMMtoccsroKORWytOYVsGYYbqut18ILWbOQfRDbyOBuzAe
IYouUztbBwLMtSFqTF2F18dW1FJ5K5QexV0qbXKn0MfwTcZ+9m6k2w9veaYIr3mQZLmr23SYkd3h
Udu8/niBXqgxxJeWimFA/oPIOIPrFjHz7qiDJ9s4u/GIae6tQXdBVbNTHOyYG0xDLhXopD6ZEi7z
HsduiqHCUrCMPmFnMY/md86ZTu5vima2SwggYefK2Ce2Tj1qnWwyHk5B/P5iNhgwCYxmwlGtkd9U
Vw6y4qt3xQ1OVXsv2Ja+ntFOZQ9EeTvK0Zd8Wx0tVcToUwmvlNvtbLfIRmbP/6jiFR1ojnNAx8J7
4SEcOuxA2Age7b3JN9TfEXzLwL72TEitjV3TgeMQyaz+isthnQPgCJ6B37+S2lpU5QVkV74wRgTL
fJ8rAOavlfwUtfFIo34oaj3N+Xd9110BPBgwi0elZTKcgjphauVxX3GfTp95DCke+fPbkv/hBEoU
opBAaLrO0S72+Hh0GP4d53K9pE3VjgphRzc1wPqI3IZdH1vQ9aLRbIUlsTsyPY9tHhCd6G1685Y7
6C341jOlNyiloev4WSn6dgiepoeJ6tOSaMcqQKgGaKOCs78ZH1dSFTO7cz7QT1ZuWUAg2gmGKrZ/
gm5DD9nPw0JGXnmYD7y1HFDAiWKbaxkMq7AIzfOQ6sERqdrZ+OP3LSlKGotw04ADjALKnbqKJwJ2
GU4shFUpw1JtRiO55NcOd8SWBXGprw/PUjVvdYWvG0AJDbBGQlZ9+ruZ0NzUW18KY7mfzIr4rLh+
nrSTAuCep+t6+s6+nOUOEwq6wH7d5zNi9ANmvBsYgk1SxzoncyY/1+OWXvKdESRqGbhgfky2MLsr
so6GH8S2BnptV4yb1epdNjBqeg7G0h9BF9G+tDx2otH5IhpbJPcznBYAKvQICNI1M+fVAOBlhzxR
x6b9Wxu1G+GXojUl68bZAbfrgHoZ9p3EGWdYjBBWQ+exDwkvOPkmvOt8J8S3zozsZvCc+9qaQgEr
orXCAdqILlWNWpnmr0xIP8XdFenMEyjVWUObxBA=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw1n;
use gw1n.components.all;

entity SPI_MASTER_Top is
port(
  I_CLK :  in std_logic;
  I_RESETN :  in std_logic;
  I_TX_EN :  in std_logic;
  I_WADDR :  in std_logic_vector(2 downto 0);
  I_WDATA :  in std_logic_vector(7 downto 0);
  I_RX_EN :  in std_logic;
  I_RADDR :  in std_logic_vector(2 downto 0);
  O_RDATA :  out std_logic_vector(7 downto 0);
  O_SPI_INT :  out std_logic;
  MISO_MASTER :  in std_logic;
  MOSI_MASTER :  out std_logic;
  SS_N_MASTER :  out std_logic_vector(3 downto 0);
  SCLK_MASTER :  out std_logic;
  MISO_SLAVE :  out std_logic;
  MOSI_SLAVE :  in std_logic;
  SS_N_SLAVE :  in std_logic;
  SCLK_SLAVE :  in std_logic);
end SPI_MASTER_Top;
architecture beh of SPI_MASTER_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
component \~spi_master.SPI_MASTER_Top\
port(
  I_CLK: in std_logic;
  I_RX_EN: in std_logic;
  MISO_MASTER: in std_logic;
  I_TX_EN: in std_logic;
  I_RESETN: in std_logic;
  I_WDATA : in std_logic_vector(7 downto 0);
  I_RADDR : in std_logic_vector(2 downto 0);
  I_WADDR : in std_logic_vector(2 downto 0);
  MOSI_MASTER: out std_logic;
  O_SPI_INT: out std_logic;
  SCLK_MASTER: out std_logic;
  O_RDATA : out std_logic_vector(7 downto 0);
  SS_N_MASTER : out std_logic_vector(3 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
u_spi_master: \~spi_master.SPI_MASTER_Top\
port map(
  I_CLK => I_CLK,
  I_RX_EN => I_RX_EN,
  MISO_MASTER => MISO_MASTER,
  I_TX_EN => I_TX_EN,
  I_RESETN => I_RESETN,
  I_WDATA(7 downto 0) => I_WDATA(7 downto 0),
  I_RADDR(2 downto 0) => I_RADDR(2 downto 0),
  I_WADDR(2 downto 0) => I_WADDR(2 downto 0),
  MOSI_MASTER => MOSI_MASTER,
  O_SPI_INT => O_SPI_INT,
  SCLK_MASTER => NN,
  O_RDATA(7 downto 0) => O_RDATA(7 downto 0),
  SS_N_MASTER(3 downto 0) => SS_N_MASTER(3 downto 0));
  SCLK_MASTER <= NN;
end beh;
